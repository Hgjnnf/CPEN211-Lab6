module cpu_tb ();